module Network (input clk, reset,
                input [63:0] inj_0, inj_1, inj_2, inj_3, inj_4, inj_5, inj_6, inj_7, inj_8, inj_9, inj_10, inj_11, inj_12, inj_13, inj_14, inj_15, 
                             inj_16, inj_17, inj_18, inj_19, inj_20, inj_21, inj_22, inj_23, inj_24, inj_25, inj_26, inj_27, inj_28, inj_29, inj_30, inj_31,
                             inj_32, inj_33, inj_34, inj_35, inj_36, inj_37, inj_38, inj_39, inj_40, inj_41, inj_42, inj_43, inj_44, inj_45, inj_46, inj_47,
                             inj_48, inj_49, inj_50, inj_51, inj_52, inj_53, inj_54, inj_55, inj_56, inj_57, inj_58, inj_59, inj_60, inj_61, inj_62, inj_63,
                output [63:0] ej_0, ej_1, ej_2, ej_3, ej_4, ej_5, ej_6, ej_7, ej_8, ej_9, ej_10, ej_11, ej_12, ej_13, ej_14, ej_15, 
                             ej_16, ej_17, ej_18, ej_19, ej_20, ej_21, ej_22, ej_23, ej_24, ej_25, ej_26, ej_27, ej_28, ej_29, ej_30, ej_31,
                             ej_32, ej_33, ej_34, ej_35, ej_36, ej_37, ej_38, ej_39, ej_40, ej_41, ej_42, ej_43, ej_44, ej_45, ej_46, ej_47,
                             ej_48, ej_49, ej_50, ej_51, ej_52, ej_53, ej_54, ej_55, ej_56, ej_57, ej_58, ej_59, ej_60, ej_61, ej_62, ej_63,
                input [63:0] push_j,
                output [63:0] write_req_j, 
                output [63:0] j_e,
                input [63:0] w_j_ack,
                output [63:0] push_j_ack);
  
 /* wire [63:0] east, west;
  wire push_w, e_state, write_req_e, w_e;
  wire push_w_ack, w_e_ack;*/
  
  wire [63:0] east [0:63];
  wire [63:0] west [0:63];
  wire [63:0] north [0:63];
  wire [63:0] south [0:63];
  
  wire E_en [0:63];
  wire W_en [0:63];
  wire N_en [0:63];
  wire S_en [0:63];
  
  wire E_req [0:63];
  wire W_req [0:63];
  wire N_req [0:63];
  wire S_req [0:63];
  
  wire E_ack [0:63];
  wire W_ack [0:63];
  wire N_ack [0:63];
  wire S_ack [0:63];
  
 /* Process_Node (input end_sim, input [2:0] X_cur, Y_cur, input [63:0] ie, iw, in, is, input clk, reset, push_e, push_w, push_n, push_s,
                     e_state, w_state, n_state, s_state, output [63:0] oe, ow, on, os, output write_req_e, write_req_w, write_req_n, write_req_s, 
                     e_e, w_e, n_e, s_e,
                     input w_e_ack, w_w_ack, w_n_ack, w_s_ack, output push_e_ack, push_w_ack, push_n_ack, push_s_ack);*/
  
  
  Process_Node p0(3'b000, 3'b000, , west[0], , south[0], clk, reset, , W_req[0], , S_req[0], E_en[0], , N_en[0], ,  east[0], , north[0], , E_req[0], , N_req[0], , , W_en[0], , S_en[0], E_ack[0], , N_ack[0], ,  , W_ack[0], , S_ack[0], inj_0, push_j[0], w_j_ack[0], write_req_j[0], j_e[0], push_j_ack[0], ej_0);
  
  Process_Node p1(3'b001, 3'b000, east[0], west[1], , south[8],  clk, reset, E_req[0], W_req[1], , S_req[8], E_en[1], W_en[0], N_en[8], , east[1], west[0], north[8], , E_req[1], W_req[0], N_req[8], , E_en[0], W_en[1], , S_en[8], E_ack[1], W_ack[0], N_ack[8], , E_ack[0], W_ack[1], , S_ack[8], inj_1, push_j[1], w_j_ack[1], write_req_j[1], j_e[1], push_j_ack[1], ej_1);
                  
  Process_Node p2(3'b010, 3'b000, east[1], west[2], , south[16],  clk, reset, E_req[1], W_req[2], , S_req[16], E_en[2], W_en[1], N_en[16], , east[2], west[1], north[16], , E_req[2], W_req[1], N_req[16], , E_en[1], W_en[2], , S_en[16], E_ack[2], W_ack[1], N_ack[16], , E_ack[1], W_ack[2], , S_ack[16], inj_2, push_j[2], w_j_ack[2], write_req_j[2], j_e[2], push_j_ack[2], ej_2);
  
  Process_Node p3(3'b011, 3'b000, east[2], west[3], , south[24],  clk, reset, E_req[2], W_req[3], , S_req[24], E_en[3], W_en[2], N_en[24], , east[3], west[2], north[24], , E_req[3], W_req[2], N_req[24], , E_en[2], W_en[3], , S_en[24], E_ack[3], W_ack[2], N_ack[24], , E_ack[2], W_ack[3], , S_ack[24], inj_3, push_j[3], w_j_ack[3], write_req_j[3], j_e[3], push_j_ack[3], ej_3);  
  
  Process_Node p4(3'b100, 3'b000, east[3], west[4], , south[32],  clk, reset, E_req[3], W_req[4], , S_req[32], E_en[4], W_en[3], N_en[32], , east[4], west[3], north[32], , E_req[4], W_req[3], N_req[32], , E_en[3], W_en[4], , S_en[32], E_ack[4], W_ack[3], N_ack[32], , E_ack[3], W_ack[4], , S_ack[32], inj_4, push_j[4], w_j_ack[4], write_req_j[4], j_e[4], push_j_ack[4], ej_4);
  
  Process_Node p5(3'b101, 3'b000, east[4], west[5], , south[40],  clk, reset, E_req[4], W_req[5], , S_req[40], E_en[5], W_en[4], N_en[40], , east[5], west[4], north[40], , E_req[5], W_req[4], N_req[40], , E_en[4], W_en[5], , S_en[40], E_ack[5], W_ack[4], N_ack[40], , E_ack[4], W_ack[5], , S_ack[40], inj_5, push_j[5], w_j_ack[5], write_req_j[5], j_e[5], push_j_ack[5], ej_5);  
  
  Process_Node p6(3'b110, 3'b000, east[5], west[6], , south[48],  clk, reset, E_req[5], W_req[6], , S_req[48], E_en[6], W_en[5], N_en[48], , east[6], west[5], north[48], , E_req[6], W_req[5], N_req[48], , E_en[5], W_en[6], , S_en[48], E_ack[6], W_ack[5], N_ack[48], , E_ack[5], W_ack[6], , S_ack[48], inj_6, push_j[6], w_j_ack[6], write_req_j[6], j_e[6], push_j_ack[6], ej_6);  
  
  Process_Node p7(3'b111, 3'b000, east[6], west[7], , south[56],  clk, reset, E_req[6], W_req[7], , S_req[56], E_en[7], W_en[6], N_en[56], , east[7], west[6], north[56], , E_req[7], W_req[6], N_req[56], , E_en[6], W_en[7], , S_en[56], E_ack[7], W_ack[6], N_ack[56], , E_ack[6], W_ack[7], , S_ack[56], inj_7, push_j[7], w_j_ack[7], write_req_j[7], j_e[7], push_j_ack[7], ej_7);  
  
  Process_Node p8(3'b000, 3'b001, , west[8], north[0], south[1],  clk, reset, , W_req[8], N_req[0], S_req[1], E_en[8], , N_en[1], S_en[0],  east[8], ,north[1] ,south[0] , E_req[8], , N_req[1], S_req[0], , W_en[8], N_en[0], S_en[1], E_ack[8], , N_ack[1], S_ack[0],  , W_ack[8], N_ack[0], S_ack[1], inj_8, push_j[8], w_j_ack[8], write_req_j[8], j_e[8], push_j_ack[8], ej_8);
  
  Process_Node p9( 3'b001, 3'b001, east[8], west[9], north[8], south[9],  clk, reset, E_req[8], W_req[9], N_req[8], S_req[9], E_en[9], W_en[8], N_en[9], S_en[8], east[9], west[8], north[9], south[8], E_req[9], W_req[8], N_req[9], S_req[8], E_en[8], W_en[9], N_en[8], S_en[9], E_ack[9], W_ack[8], N_ack[9], S_ack[8], E_ack[8], W_ack[9], N_ack[8], S_ack[9], inj_9, push_j[9], w_j_ack[9], write_req_j[9], j_e[9], push_j_ack[9], ej_9);
                  
  Process_Node p10( 3'b010, 3'b001, east[9], west[10], north[16], south[17], clk, reset, E_req[9], W_req[10], N_req[16], S_req[17], E_en[10], W_en[9], N_en[17], S_en[16], east[10], west[9], north[17], south[16], E_req[10], W_req[9], N_req[17], S_req[16], E_en[9], W_en[10], N_en[16], S_en[17], E_ack[10], W_ack[9], N_ack[17], S_ack[16], E_ack[9], W_ack[10], N_ack[16], S_ack[17], inj_10, push_j[10], w_j_ack[10], write_req_j[10], j_e[10], push_j_ack[10], ej_10);
  
  Process_Node p11( 3'b011, 3'b001, east[10], west[11], north[24], south[25], clk, reset, E_req[10], W_req[11], N_req[24], S_req[25], E_en[11], W_en[10], N_en[25], S_en[24], east[11], west[10], north[25], south[24], E_req[11], W_req[10], N_req[25], S_req[24], E_en[10], W_en[11], N_en[24], S_en[25], E_ack[11], W_ack[10], N_ack[25], S_ack[24], E_ack[10], W_ack[11], N_ack[24], S_ack[25], inj_11, push_j[11], w_j_ack[11], write_req_j[11], j_e[11], push_j_ack[11], ej_11);  
  
  Process_Node p12( 3'b100, 3'b001, east[11], west[12], north[32], south[33], clk, reset, E_req[11], W_req[12], N_req[32], S_req[33], E_en[12], W_en[11], N_en[33], S_en[32], east[12], west[11], north[33], south[32], E_req[12], W_req[11], N_req[33], S_req[32], E_en[11], W_en[12], N_en[32], S_en[33], E_ack[12], W_ack[11], N_ack[33], S_ack[32], E_ack[11], W_ack[12], N_ack[32], S_ack[33], inj_12, push_j[12], w_j_ack[12], write_req_j[12], j_e[12], push_j_ack[12], ej_12);
  
  Process_Node p13( 3'b101, 3'b001, east[12], west[13], north[40], south[41], clk, reset, E_req[12], W_req[13], N_req[40], S_req[41], E_en[13], W_en[12], N_en[41], S_en[40], east[13], west[12], north[41], south[40], E_req[13], W_req[12], N_req[41], S_req[40], E_en[12], W_en[13], N_en[40], S_en[41], E_ack[13], W_ack[12], N_ack[41], S_ack[40], E_ack[12], W_ack[13], N_ack[40], S_ack[41], inj_13, push_j[13], w_j_ack[13], write_req_j[13], j_e[13], push_j_ack[13], ej_13);  
  
  Process_Node p14( 3'b110, 3'b001, east[13], west[14], north[48], south[49], clk, reset, E_req[13], W_req[14], N_req[48], S_req[49], E_en[14], W_en[13], N_en[49], S_en[48], east[14], west[13], north[49], south[48], E_req[14], W_req[13], N_req[49], S_req[48], E_en[13], W_en[14], N_en[48], S_en[49], E_ack[14], W_ack[13], N_ack[49], S_ack[48], E_ack[13], W_ack[14], N_ack[48], S_ack[49], inj_14, push_j[14], w_j_ack[14], write_req_j[14], j_e[14], push_j_ack[14], ej_14);  
  
  Process_Node p15( 3'b111, 3'b001, east[14], west[15], north[56], south[57], clk, reset, E_req[14], W_req[15], N_req[56], S_req[57], E_en[15], W_en[14], N_en[57], S_en[56], east[15], west[14], north[57], south[56], E_req[15], W_req[14], N_req[57], S_req[56], E_en[14], W_en[15], N_en[56], S_en[57], E_ack[15], W_ack[14], N_ack[57], S_ack[56], E_ack[14], W_ack[15], N_ack[56], S_ack[57], inj_15, push_j[15], w_j_ack[15], write_req_j[15], j_e[15], push_j_ack[15], ej_15);  
  
  Process_Node p16( 3'b000, 3'b010, , west[16], north[1], south[2],  clk, reset, , W_req[16], N_req[1], S_req[2], E_en[16], , N_en[2], S_en[1],  east[16], , north[2], south[1], E_req[16], , N_req[2], S_req[1], , W_en[16], N_en[1], S_en[2], E_ack[16], , N_ack[2], S_ack[1],  , W_ack[16], N_ack[1], S_ack[2], inj_16, push_j[16], w_j_ack[16], write_req_j[16], j_e[16], push_j_ack[16], ej_16);
  
  Process_Node p17( 3'b001, 3'b010, east[16], west[17], north[9], south[10],  clk, reset, E_req[16], W_req[17], N_req[9], S_req[10], E_en[17], W_en[16], N_en[10], S_en[9], east[17], west[16], north[10], south[9], E_req[17], W_req[16], N_req[10], S_req[9], E_en[16], W_en[17], N_en[9], S_en[10], E_ack[17], W_ack[16], N_ack[10], S_ack[9], E_ack[16], W_ack[17], N_ack[9], S_ack[10], inj_17, push_j[17], w_j_ack[17], write_req_j[17], j_e[17], push_j_ack[17], ej_17);
                  
  Process_Node p18( 3'b010, 3'b010, east[17], west[18], north[17], south[18], clk, reset, E_req[17], W_req[18], N_req[17], S_req[18], E_en[18], W_en[17], N_en[18], S_en[17], east[18], west[17], north[18], south[17], E_req[18], W_req[17], N_req[18], S_req[17], E_en[17], W_en[18], N_en[17], S_en[18], E_ack[18], W_ack[17], N_ack[18], S_ack[17], E_ack[17], W_ack[18], N_ack[17], S_ack[18], inj_18, push_j[18], w_j_ack[18], write_req_j[18], j_e[18], push_j_ack[18], ej_18);
  
  Process_Node p19( 3'b011, 3'b010, east[18], west[19], north[25], south[26], clk, reset, E_req[18], W_req[19], N_req[25], S_req[26], E_en[19], W_en[18], N_en[26], S_en[25], east[19], west[18], north[26], south[25], E_req[19], W_req[18], N_req[26], S_req[25], E_en[18], W_en[19], N_en[25], S_en[26], E_ack[19], W_ack[18], N_ack[26], S_ack[25], E_ack[18], W_ack[19], N_ack[25], S_ack[26], inj_19, push_j[19], w_j_ack[19], write_req_j[19], j_e[19], push_j_ack[19], ej_19);  
  
  Process_Node p20( 3'b100, 3'b010, east[19], west[20], north[33], south[34], clk, reset, E_req[19], W_req[20], N_req[33], S_req[34], E_en[20], W_en[19], N_en[34], S_en[33], east[20], west[19], north[34], south[33], E_req[20], W_req[19], N_req[34], S_req[33], E_en[19], W_en[20], N_en[33], S_en[34], E_ack[20], W_ack[19], N_ack[34], S_ack[33], E_ack[19], W_ack[20], N_ack[33], S_ack[34], inj_20, push_j[20], w_j_ack[20], write_req_j[20], j_e[20], push_j_ack[20], ej_20);
  
  Process_Node p21( 3'b101, 3'b010, east[20], west[21], north[41], south[42], clk, reset, E_req[20], W_req[21], N_req[41], S_req[42], E_en[21], W_en[20], N_en[42], S_en[41], east[21], west[20], north[42], south[41], E_req[21], W_req[20], N_req[42], S_req[41], E_en[20], W_en[21], N_en[41], S_en[42], E_ack[21], W_ack[20], N_ack[42], S_ack[41], E_ack[20], W_ack[21], N_ack[41], S_ack[42], inj_21, push_j[21], w_j_ack[21], write_req_j[21], j_e[21], push_j_ack[21], ej_21);  
  
  Process_Node p22( 3'b110, 3'b010, east[21], west[22], north[49], south[50], clk, reset, E_req[21], W_req[22], N_req[49], S_req[50], E_en[22], W_en[21], N_en[50], S_en[49], east[22], west[21], north[50], south[49], E_req[22], W_req[21], N_req[50], S_req[49], E_en[21], W_en[22], N_en[49], S_en[50], E_ack[22], W_ack[21], N_ack[50], S_ack[49], E_ack[21], W_ack[22], N_ack[49], S_ack[50], inj_22, push_j[22], w_j_ack[22], write_req_j[22], j_e[22], push_j_ack[22], ej_22);  
  
  Process_Node p23( 3'b111, 3'b010, east[22], west[23], north[57], south[58], clk, reset, E_req[22], W_req[23], N_req[57], S_req[58], E_en[23], W_en[22], N_en[58], S_en[57], east[23], west[22], north[58], south[57], E_req[23], W_req[22], N_req[58], S_req[57], E_en[22], W_en[23], N_en[57], S_en[58], E_ack[23], W_ack[22], N_ack[58], S_ack[57], E_ack[22], W_ack[23], N_ack[57], S_ack[58], inj_23, push_j[23], w_j_ack[23], write_req_j[23], j_e[23], push_j_ack[23], ej_23);  
  
  Process_Node p24( 3'b000, 3'b011, , west[24], north[2], south[3],  clk, reset, , W_req[24], N_req[2], S_req[3], E_en[24], , N_en[3], S_en[2], east[24], , north[3], south[2], E_req[24], , N_req[3], S_req[2], , W_en[24], N_en[2], S_en[3], E_ack[24], , N_ack[3], S_ack[2],  , W_ack[24], N_ack[2], S_ack[3], inj_24, push_j[24], w_j_ack[24], write_req_j[24], j_e[24], push_j_ack[24], ej_24);
  
  Process_Node p25( 3'b001, 3'b011, east[24], west[25], north[10], south[11],  clk, reset, E_req[24], W_req[25], N_req[10], S_req[11], E_en[25], W_en[24], N_en[11], S_en[10], east[25], west[24], north[11], south[10], E_req[25], W_req[24], N_req[11], S_req[10], E_en[24], W_en[25], N_en[10], S_en[11], E_ack[25], W_ack[24], N_ack[11], S_ack[10], E_ack[24], W_ack[25], N_ack[10], S_ack[11], inj_25, push_j[25], w_j_ack[25], write_req_j[25], j_e[25], push_j_ack[25], ej_25);
                  
  Process_Node p26( 3'b010, 3'b011, east[25], west[26], north[18], south[19], clk, reset, E_req[25], W_req[26], N_req[18], S_req[19], E_en[26], W_en[25], N_en[19], S_en[18], east[26], west[25], north[19], south[18], E_req[26], W_req[25], N_req[19], S_req[18], E_en[25], W_en[26], N_en[18], S_en[19], E_ack[26], W_ack[25], N_ack[19], S_ack[18], E_ack[25], W_ack[26], N_ack[18], S_ack[19], inj_26, push_j[26], w_j_ack[26], write_req_j[26], j_e[26], push_j_ack[26], ej_26);
  
  Process_Node p27( 3'b011, 3'b011, east[26], west[27], north[26], south[27], clk, reset, E_req[26], W_req[27], N_req[26], S_req[27], E_en[27], W_en[26], N_en[27], S_en[26], east[27], west[26], north[27], south[26], E_req[27], W_req[26], N_req[27], S_req[26], E_en[26], W_en[27], N_en[26], S_en[27], E_ack[27], W_ack[26], N_ack[27], S_ack[26], E_ack[26], W_ack[27], N_ack[26], S_ack[27], inj_27, push_j[27], w_j_ack[27], write_req_j[27], j_e[27], push_j_ack[27], ej_27);  
  
  Process_Node p28( 3'b100, 3'b011, east[27], west[28], north[34], south[35], clk, reset, E_req[27], W_req[28], N_req[34], S_req[35], E_en[28], W_en[27], N_en[35], S_en[34], east[28], west[27], north[35], south[34], E_req[28], W_req[27], N_req[35], S_req[34], E_en[27], W_en[28], N_en[34], S_en[35], E_ack[28], W_ack[27], N_ack[35], S_ack[34], E_ack[27], W_ack[28], N_ack[34], S_ack[35], inj_28, push_j[28], w_j_ack[28], write_req_j[28], j_e[28], push_j_ack[28], ej_28);
  
  Process_Node p29( 3'b101, 3'b011, east[28], west[29], north[42], south[43], clk, reset, E_req[28], W_req[29], N_req[42], S_req[43], E_en[29], W_en[28], N_en[43], S_en[42], east[29], west[28], north[43], south[42], E_req[29], W_req[28], N_req[43], S_req[42], E_en[28], W_en[29], N_en[42], S_en[43], E_ack[29], W_ack[28], N_ack[43], S_ack[42], E_ack[28], W_ack[29], N_ack[42], S_ack[43], inj_29, push_j[29], w_j_ack[29], write_req_j[29], j_e[29], push_j_ack[29], ej_29);  
  
  Process_Node p30( 3'b110, 3'b011, east[29], west[30], north[50], south[51], clk, reset, E_req[29], W_req[30], N_req[50], S_req[51], E_en[30], W_en[29], N_en[51], S_en[50], east[30], west[29], north[51], south[50], E_req[30], W_req[29], N_req[51], S_req[50], E_en[29], W_en[30], N_en[50], S_en[51], E_ack[30], W_ack[29], N_ack[51], S_ack[50], E_ack[29], W_ack[30], N_ack[50], S_ack[51], inj_30, push_j[30], w_j_ack[30], write_req_j[30], j_e[30], push_j_ack[30], ej_30);  
  
  Process_Node p31( 3'b111, 3'b011, east[30], west[31], north[58], south[59], clk, reset, E_req[30], W_req[31], N_req[58], S_req[59], E_en[31], W_en[30], N_en[59], S_en[58], east[31], west[30], north[59], south[58], E_req[31], W_req[30], N_req[59], S_req[58], E_en[30], W_en[31], N_en[58], S_en[59], E_ack[31], W_ack[30], N_ack[59], S_ack[58], E_ack[30], W_ack[31], N_ack[58], S_ack[59], inj_31, push_j[31], w_j_ack[31], write_req_j[31], j_e[31], push_j_ack[31], ej_31);  
  
  Process_Node p32( 3'b000, 3'b100, , west[32], north[3], south[4],  clk, reset, , W_req[32], N_req[3], S_req[4], E_en[32], , N_en[4], S_en[3],  east[32], , north[4], south[3], E_req[32], , N_req[4], S_req[3], , W_en[32], N_en[3], S_en[4], E_ack[32], , N_ack[4], S_ack[3],  , W_ack[32], N_ack[3], S_ack[4], inj_32, push_j[32], w_j_ack[32], write_req_j[32], j_e[32], push_j_ack[32], ej_32);
  
  Process_Node p33( 3'b001, 3'b100, east[32], west[33], north[11], south[12],  clk, reset, E_req[32], W_req[33], N_req[11], S_req[12], E_en[33], W_en[32], N_en[12], S_en[11], east[33], west[32], north[12], south[11], E_req[33], W_req[32], N_req[12], S_req[11], E_en[32], W_en[33], N_en[11], S_en[12], E_ack[33], W_ack[32], N_ack[12], S_ack[11], E_ack[32], W_ack[33], N_ack[11], S_ack[12], inj_33, push_j[33], w_j_ack[33], write_req_j[33], j_e[33], push_j_ack[33], ej_33);
                  
  Process_Node p34( 3'b010, 3'b100, east[33], west[34], north[19], south[20], clk, reset, E_req[33], W_req[34], N_req[19], S_req[20], E_en[34], W_en[33], N_en[20], S_en[19], east[34], west[33], north[20], south[19], E_req[34], W_req[33], N_req[20], S_req[19], E_en[33], W_en[34], N_en[19], S_en[20], E_ack[34], W_ack[33], N_ack[20], S_ack[19], E_ack[33], W_ack[34], N_ack[19], S_ack[20], inj_34, push_j[34], w_j_ack[34], write_req_j[34], j_e[34], push_j_ack[34], ej_34);
  
  Process_Node p35( 3'b011, 3'b100, east[34], west[35], north[27], south[28], clk, reset, E_req[34], W_req[35], N_req[27], S_req[28], E_en[35], W_en[34], N_en[28], S_en[27], east[35], west[34], north[28], south[27], E_req[35], W_req[34], N_req[28], S_req[27], E_en[34], W_en[35], N_en[27], S_en[28], E_ack[35], W_ack[34], N_ack[28], S_ack[27], E_ack[34], W_ack[35], N_ack[27], S_ack[28], inj_35, push_j[35], w_j_ack[35], write_req_j[35], j_e[35], push_j_ack[35], ej_35);  
  
  Process_Node p36( 3'b100, 3'b100, east[35], west[36], north[35], south[36], clk, reset, E_req[35], W_req[36], N_req[35], S_req[36], E_en[36], W_en[35], N_en[36], S_en[35], east[36], west[35], north[36], south[35], E_req[36], W_req[35], N_req[36], S_req[35], E_en[35], W_en[36], N_en[35], S_en[36], E_ack[36], W_ack[35], N_ack[36], S_ack[35], E_ack[35], W_ack[36], N_ack[35], S_ack[36], inj_36, push_j[36], w_j_ack[36], write_req_j[36], j_e[36], push_j_ack[36], ej_36);
  
  Process_Node p37( 3'b101, 3'b100, east[36], west[37], north[43], south[44], clk, reset, E_req[36], W_req[37], N_req[43], S_req[44], E_en[37], W_en[36], N_en[44], S_en[43], east[37], west[36], north[44], south[43], E_req[37], W_req[36], N_req[44], S_req[43], E_en[36], W_en[37], N_en[43], S_en[44], E_ack[37], W_ack[36], N_ack[44], S_ack[43], E_ack[36], W_ack[37], N_ack[43], S_ack[44], inj_37, push_j[37], w_j_ack[37], write_req_j[37], j_e[37], push_j_ack[37], ej_37);  
  
  Process_Node p38( 3'b110, 3'b100, east[37], west[38], north[51], south[52], clk, reset, E_req[37], W_req[38], N_req[51], S_req[52], E_en[38], W_en[37], N_en[52], S_en[51], east[38], west[37], north[52], south[51], E_req[38], W_req[37], N_req[52], S_req[51], E_en[37], W_en[38], N_en[51], S_en[52], E_ack[38], W_ack[37], N_ack[52], S_ack[51], E_ack[37], W_ack[38], N_ack[51], S_ack[52], inj_38, push_j[38], w_j_ack[38], write_req_j[38], j_e[38], push_j_ack[38], ej_38);  
  
  Process_Node p39( 3'b111, 3'b100, east[38], west[39], north[59], south[60], clk, reset, E_req[38], W_req[39], N_req[59], S_req[60], E_en[39], W_en[38], N_en[60], S_en[59], east[39], west[38], north[60], south[59], E_req[39], W_req[38], N_req[60], S_req[59], E_en[38], W_en[39], N_en[59], S_en[60], E_ack[39], W_ack[38], N_ack[60], S_ack[59], E_ack[38], W_ack[39], N_ack[59], S_ack[60], inj_39, push_j[39], w_j_ack[39], write_req_j[39], j_e[39], push_j_ack[39], ej_39);  
  
  Process_Node p40( 3'b000, 3'b101, , west[40], north[4], south[5],  clk, reset, , W_req[40], N_req[4], S_req[5], E_en[40], , N_en[5], S_en[4],  east[40], , north[5], south[4], E_req[40], , N_req[5], S_req[4], , W_en[40], N_en[4], S_en[5], E_ack[40], , N_ack[5], S_ack[4],  , W_ack[40], N_ack[4], S_ack[5], inj_40, push_j[40], w_j_ack[40], write_req_j[40], j_e[40], push_j_ack[40], ej_40);
  
  Process_Node p41( 3'b001, 3'b101, east[40], west[41], north[12], south[13],  clk, reset, E_req[40], W_req[41], N_req[12], S_req[13], E_en[41], W_en[40], N_en[13], S_en[12], east[41], west[40], north[13], south[12], E_req[41], W_req[40], N_req[13], S_req[12], E_en[40], W_en[41], N_en[12], S_en[13], E_ack[41], W_ack[40], N_ack[13], S_ack[12], E_ack[40], W_ack[41], N_ack[12], S_ack[13], inj_41, push_j[41], w_j_ack[41], write_req_j[41], j_e[41], push_j_ack[41], ej_41);
                  
  Process_Node p42( 3'b010, 3'b101, east[41], west[42], north[20], south[21], clk, reset, E_req[41], W_req[42], N_req[20], S_req[21], E_en[42], W_en[41], N_en[21], S_en[20], east[42], west[41], north[21], south[20], E_req[42], W_req[41], N_req[21], S_req[20], E_en[41], W_en[42], N_en[20], S_en[21], E_ack[42], W_ack[41], N_ack[21], S_ack[20], E_ack[41], W_ack[42], N_ack[20], S_ack[21], inj_42, push_j[42], w_j_ack[42], write_req_j[42], j_e[42], push_j_ack[42], ej_42);
  
  Process_Node p43( 3'b011, 3'b101, east[42], west[43], north[28], south[29], clk, reset, E_req[42], W_req[43], N_req[28], S_req[29], E_en[43], W_en[42], N_en[29], S_en[28], east[43], west[42], north[29], south[28], E_req[43], W_req[42], N_req[29], S_req[28], E_en[42], W_en[43], N_en[28], S_en[29], E_ack[43], W_ack[42], N_ack[29], S_ack[28], E_ack[42], W_ack[43], N_ack[28], S_ack[29], inj_43, push_j[43], w_j_ack[43], write_req_j[43], j_e[43], push_j_ack[43], ej_43);  
  
  Process_Node p44( 3'b100, 3'b101, east[43], west[44], north[36], south[37], clk, reset, E_req[43], W_req[44], N_req[36], S_req[37], E_en[44], W_en[43], N_en[37], S_en[36], east[44], west[43], north[37], south[36], E_req[44], W_req[43], N_req[37], S_req[36], E_en[43], W_en[44], N_en[36], S_en[37], E_ack[44], W_ack[43], N_ack[37], S_ack[36], E_ack[43], W_ack[44], N_ack[36], S_ack[37], inj_44, push_j[44], w_j_ack[44], write_req_j[44], j_e[44], push_j_ack[44], ej_44);
  
  Process_Node p45( 3'b101, 3'b101, east[44], west[45], north[44], south[45], clk, reset, E_req[44], W_req[45], N_req[44], S_req[45], E_en[45], W_en[44], N_en[45], S_en[44], east[45], west[44], north[45], south[44], E_req[45], W_req[44], N_req[45], S_req[44], E_en[44], W_en[45], N_en[44], S_en[45], E_ack[45], W_ack[44], N_ack[45], S_ack[44], E_ack[44], W_ack[45], N_ack[44], S_ack[45], inj_45, push_j[45], w_j_ack[45], write_req_j[45], j_e[45], push_j_ack[45], ej_45);  
  
  Process_Node p46( 3'b110, 3'b101, east[45], west[46], north[52], south[53], clk, reset, E_req[45], W_req[46], N_req[52], S_req[53], E_en[46], W_en[45], N_en[53], S_en[52], east[46], west[45], north[53], south[52], E_req[46], W_req[45], N_req[53], S_req[52], E_en[45], W_en[46], N_en[52], S_en[53], E_ack[46], W_ack[45], N_ack[53], S_ack[52], E_ack[45], W_ack[46], N_ack[52], S_ack[53], inj_46, push_j[46], w_j_ack[46], write_req_j[46], j_e[46], push_j_ack[46], ej_46);  
  
  Process_Node p47( 3'b111, 3'b101, east[46], west[47], north[60], south[61], clk, reset, E_req[46], W_req[47], N_req[60], S_req[61], E_en[47], W_en[46], N_en[61], S_en[60], east[47], west[46], north[61], south[60], E_req[47], W_req[46], N_req[61], S_req[60], E_en[46], W_en[47], N_en[60], S_en[61], E_ack[47], W_ack[46], N_ack[61], S_ack[60], E_ack[46], W_ack[47], N_ack[60], S_ack[61], inj_47, push_j[47], w_j_ack[47], write_req_j[47], j_e[47], push_j_ack[47], ej_47);  
  
  Process_Node p48( 3'b000, 3'b110, , west[48], north[5], south[6],  clk, reset, , W_req[48], N_req[5], S_req[6], E_en[48], , N_en[6], S_en[5],  east[48], , north[6], south[5], E_req[48], , N_req[6], S_req[5], , W_en[48], N_en[5], S_en[6], E_ack[48], , N_ack[6], S_ack[5],  , W_ack[48], N_ack[5], S_ack[6], inj_48, push_j[48], w_j_ack[48], write_req_j[48], j_e[48], push_j_ack[48], ej_48);
  
  Process_Node p49( 3'b001, 3'b110, east[48], west[49], north[13], south[14],  clk, reset, E_req[48], W_req[49], N_req[13], S_req[14], E_en[49], W_en[48], N_en[14], S_en[13], east[49], west[48], north[14], south[13], E_req[49], W_req[48], N_req[14], S_req[13], E_en[48], W_en[49], N_en[13], S_en[14], E_ack[49], W_ack[48], N_ack[14], S_ack[13], E_ack[48], W_ack[49], N_ack[13], S_ack[14], inj_49, push_j[49], w_j_ack[49], write_req_j[49], j_e[49], push_j_ack[49], ej_49);
                  
  Process_Node p50( 3'b010, 3'b110, east[49], west[50], north[21], south[22], clk, reset, E_req[49], W_req[50], N_req[21], S_req[22], E_en[50], W_en[49], N_en[22], S_en[21], east[50], west[49], north[22], south[21], E_req[50], W_req[49], N_req[22], S_req[21], E_en[49], W_en[50], N_en[21], S_en[22], E_ack[50], W_ack[49], N_ack[22], S_ack[21], E_ack[49], W_ack[50], N_ack[21], S_ack[22], inj_50, push_j[50], w_j_ack[50], write_req_j[50], j_e[50], push_j_ack[50], ej_50);
  
  Process_Node p51( 3'b011, 3'b110, east[50], west[51], north[29], south[30], clk, reset, E_req[50], W_req[51], N_req[29], S_req[30], E_en[51], W_en[50], N_en[30], S_en[29], east[51], west[50], north[30], south[29], E_req[51], W_req[50], N_req[30], S_req[29], E_en[50], W_en[51], N_en[29], S_en[30], E_ack[51], W_ack[50], N_ack[30], S_ack[29], E_ack[50], W_ack[51], N_ack[29], S_ack[30], inj_51, push_j[51], w_j_ack[51], write_req_j[51], j_e[51], push_j_ack[51], ej_51);  
  
  Process_Node p52( 3'b100, 3'b110, east[51], west[52], north[37], south[38], clk, reset, E_req[51], W_req[52], N_req[37], S_req[38], E_en[52], W_en[51], N_en[38], S_en[37], east[52], west[51], north[38], south[37], E_req[52], W_req[51], N_req[38], S_req[37], E_en[51], W_en[52], N_en[37], S_en[38], E_ack[52], W_ack[51], N_ack[38], S_ack[37], E_ack[51], W_ack[52], N_ack[37], S_ack[38], inj_52, push_j[52], w_j_ack[52], write_req_j[52], j_e[52], push_j_ack[52], ej_52);
  
  Process_Node p53( 3'b101, 3'b110, east[52], west[53], north[45], south[46], clk, reset, E_req[52], W_req[53], N_req[45], S_req[46], E_en[53], W_en[52], N_en[46], S_en[45], east[53], west[52], north[46], south[45], E_req[53], W_req[52], N_req[46], S_req[45], E_en[52], W_en[53], N_en[45], S_en[46], E_ack[53], W_ack[52], N_ack[46], S_ack[45], E_ack[52], W_ack[53], N_ack[45], S_ack[46], inj_53, push_j[53], w_j_ack[53], write_req_j[53], j_e[53], push_j_ack[53], ej_53);  
  
  Process_Node p54( 3'b110, 3'b110, east[53], west[54], north[53], south[54], clk, reset, E_req[53], W_req[54], N_req[53], S_req[54], E_en[54], W_en[53], N_en[54], S_en[53], east[54], west[53], north[54], south[53], E_req[54], W_req[53], N_req[54], S_req[53], E_en[53], W_en[54], N_en[53], S_en[54], E_ack[54], W_ack[53], N_ack[54], S_ack[53], E_ack[53], W_ack[54], N_ack[53], S_ack[54], inj_54, push_j[54], w_j_ack[54], write_req_j[54], j_e[54], push_j_ack[54], ej_54);  
  
  Process_Node p55( 3'b111, 3'b110, east[54], west[55], north[61], south[62], clk, reset, E_req[54], W_req[55], N_req[61], S_req[62], E_en[55], W_en[54], N_en[62], S_en[61], east[55], west[54], north[62], south[61], E_req[55], W_req[54], N_req[62], S_req[61], E_en[54], W_en[55], N_en[61], S_en[62], E_ack[55], W_ack[54], N_ack[62], S_ack[61], E_ack[54], W_ack[55], N_ack[61], S_ack[62], inj_55, push_j[55], w_j_ack[55], write_req_j[55], j_e[55], push_j_ack[55], ej_55);  
  
  Process_Node p56( 3'b000, 3'b111, , west[56], north[6], south[7],  clk, reset, , W_req[56], N_req[6], S_req[7], E_en[56], , N_en[7], S_en[6],  east[56], , north[7], south[6], E_req[56], , N_req[7], S_req[6], , W_en[56], N_en[6], S_en[7], E_ack[56], , N_ack[7], S_ack[6],  , W_ack[56], N_ack[6], S_ack[7], inj_56, push_j[56], w_j_ack[56], write_req_j[56], j_e[56], push_j_ack[56], ej_56);
  
  Process_Node p57( 3'b001, 3'b111, east[56], west[57], north[14], south[15],  clk, reset, E_req[56], W_req[57], N_req[14], S_req[15], E_en[57], W_en[56], N_en[15], S_en[14], east[57], west[56], north[15], south[14], E_req[57], W_req[56], N_req[15], S_req[14], E_en[56], W_en[57], N_en[14], S_en[15], E_ack[57], W_ack[56], N_ack[15], S_ack[14], E_ack[56], W_ack[57], N_ack[14], S_ack[15], inj_57, push_j[57], w_j_ack[57], write_req_j[57], j_e[57], push_j_ack[57], ej_57);
                  
  Process_Node p58( 3'b010, 3'b111, east[57], west[58], north[22], south[23], clk, reset, E_req[57], W_req[58], N_req[22], S_req[23], E_en[58], W_en[57], N_en[23], S_en[22], east[58], west[57], north[23], south[22], E_req[58], W_req[57], N_req[23], S_req[22], E_en[57], W_en[58], N_en[22], S_en[23], E_ack[58], W_ack[57], N_ack[23], S_ack[22], E_ack[57], W_ack[58], N_ack[22], S_ack[23], inj_58, push_j[58], w_j_ack[58], write_req_j[58], j_e[58], push_j_ack[58], ej_58);
  
  Process_Node p59( 3'b011, 3'b111, east[58], west[59], north[30], south[31], clk, reset, E_req[58], W_req[59], N_req[30], S_req[31], E_en[59], W_en[58], N_en[31], S_en[30], east[59], west[58], north[31], south[30], E_req[59], W_req[58], N_req[31], S_req[30], E_en[58], W_en[59], N_en[30], S_en[31], E_ack[59], W_ack[58], N_ack[31], S_ack[30], E_ack[58], W_ack[59], N_ack[30], S_ack[31], inj_59, push_j[59], w_j_ack[59], write_req_j[59], j_e[59], push_j_ack[59], ej_59);  
  
  Process_Node p60( 3'b100, 3'b111, east[59], west[60], north[38], south[39], clk, reset, E_req[59], W_req[60], N_req[38], S_req[39], E_en[60], W_en[59], N_en[39], S_en[38], east[60], west[59], north[39], south[38], E_req[60], W_req[59], N_req[39], S_req[38], E_en[59], W_en[60], N_en[38], S_en[39], E_ack[60], W_ack[59], N_ack[39], S_ack[38], E_ack[59], W_ack[60], N_ack[38], S_ack[39], inj_60, push_j[60], w_j_ack[60], write_req_j[60], j_e[60], push_j_ack[60], ej_60);
  
  Process_Node p61( 3'b101, 3'b111, east[60], west[61], north[46], south[47], clk, reset, E_req[60], W_req[61], N_req[46], S_req[47], E_en[61], W_en[60], N_en[47], S_en[46], east[61], west[60], north[47], south[46], E_req[61], W_req[60], N_req[47], S_req[46], E_en[60], W_en[61], N_en[46], S_en[47], E_ack[61], W_ack[60], N_ack[47], S_ack[46], E_ack[60], W_ack[61], N_ack[46], S_ack[47], inj_61, push_j[61], w_j_ack[61], write_req_j[61], j_e[61], push_j_ack[61], ej_61);  
  
  Process_Node p62( 3'b110, 3'b111, east[61], west[62], north[54], south[55], clk, reset, E_req[61], W_req[62], N_req[54], S_req[55], E_en[62], W_en[61], N_en[55], S_en[54], east[62], west[61], north[55], south[54], E_req[62], W_req[61], N_req[55], S_req[54], E_en[61], W_en[62], N_en[54], S_en[55], E_ack[62], W_ack[61], N_ack[55], S_ack[54], E_ack[61], W_ack[62], N_ack[54], S_ack[55], inj_62, push_j[62], w_j_ack[62], write_req_j[62], j_e[62], push_j_ack[62], ej_62);  
  
  Process_Node p63( 3'b111, 3'b111, east[62], west[63], north[62], south[63], clk, reset, E_req[62], W_req[63], N_req[62], S_req[63], E_en[63], W_en[62], N_en[63], S_en[62], east[63], west[62], north[63], south[62], E_req[63], W_req[62], N_req[63], S_req[62], E_en[62], W_en[63], N_en[62], S_en[63], E_ack[63], W_ack[62], N_ack[63], S_ack[62], E_ack[62], W_ack[63], N_ack[62], S_ack[63], inj_63, push_j[63], w_j_ack[63], write_req_j[63], j_e[63], push_j_ack[63], ej_63);  
  
  
endmodule
